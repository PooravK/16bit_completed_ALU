module arith_top();
endmodule