module alu_top();

endmodule