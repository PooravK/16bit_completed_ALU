parameter ALU_ADD = 5'b00000;
parameter ALU_SUB = 5'b00001;
parameter ALU_MUL = 5'b00010;
parameter ALU_DIV = 5'b00011;

parameter ALU_AND = 5'b01000;
parameter ALU_OR  = 5'b01001;
parameter ALU_XOR = 5'b01010;
parameter ALU_NOT = 5'b01011;
parameter ALU_NAND= 5'b01100;
parameter ALU_NOR = 5'b01101;
parameter ALU_XNOR= 5'b01110;

parameter ALU_UNSIGNED_GT = 5'b10000;
parameter ALU_SIGNED_GT   = 5'b10001;
parameter ALU_UNSIGNED_LT = 5'b10010;
parameter ALU_SIGNED_LT   = 5'b10011;
parameter ALU_UNSIGNED_ET = 5'b10100;
parameter ALU_SIGNED_ET   = 5'b10101;

parameter ALU_LSL = 5'b11000;
parameter ALU_LSR = 5'b11001;
parameter ALU_ASL = 5'b11010;
parameter ALU_ASR = 5'b11011;
parameter ALU_RL  = 5'b11100;
parameter ALU_RR  = 5'b11101;