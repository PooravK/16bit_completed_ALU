module signed_mult(
    );
endmodule