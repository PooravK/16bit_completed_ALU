module signed_mult(
    input [15:0]in0, in1,
    output [31:0]s_prod
    );
endmodule